--Mitchell Irvin
--Small8
--Section: 1525
--Small8 Datapath TB

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity datapath_tb is
end datapath_tb;

architecture tb of datapath_tb is
begin


end tb; 